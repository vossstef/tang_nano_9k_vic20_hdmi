--Copyright (C)2014-2022 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.09 Education
--Part Number: GW1NR-LV9QN88PC6/I5
--Device: GW1NR-9C
--Created Time: Mon Jan 16 12:50:26 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_char is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(11 downto 0)
    );
end Gowin_pROM_char;

architecture Behavioral of Gowin_pROM_char is

    signal prom_inst_0_dout_w: std_logic_vector(27 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(27 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(11 downto 0) & gw_gnd & gw_gnd;
    dout(3 downto 0) <= prom_inst_0_DO_o(3 downto 0) ;
    prom_inst_0_dout_w(27 downto 0) <= prom_inst_0_DO_o(31 downto 4) ;
    prom_inst_1_AD_i <= ad(11 downto 0) & gw_gnd & gw_gnd;
    dout(7 downto 4) <= prom_inst_1_DO_o(3 downto 0) ;
    prom_inst_1_dout_w(27 downto 0) <= prom_inst_1_DO_o(31 downto 4) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 4,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0C22E02C0000800E0E00800E084222480C20002C0C22C22C0222E2480E0C6A2C",
            INIT_RAM_01 => X"084222480226A2220222AA620E000000024808420844444E0C88888C0222E222",
            INIT_RAM_02 => X"026AA222088442220C2222220888888E0C22C02C0248C22C0A4A22480000C22C",
            INIT_RAM_03 => X"000F00008888AC800C44444C0E00C00C0C00000C0E00842E0888C22202248422",
            INIT_RAM_04 => X"000000840A4A08800660842008CAC8E8044E4E44000004440800888800000000",
            INIT_RAM_05 => X"00008420088000000000E000088000000088E88008ACECA80008880004800084",
            INIT_RAM_06 => X"0000842E0C22C00C0842480E044E44C40C22C22C0E00C22C0E8888880C22A62C",
            INIT_RAM_07 => X"0000C22C008C6C80000E0E000E80008E08800800008008000842E22C0C22C22C",
            INIT_RAM_08 => X"0000000000F00000000000F000000F000000F000000000000ECFFEC8000F0000",
            INIT_RAM_09 => X"0000000F0000842112480000F000000000000888000348888800000044444444",
            INIT_RAM_0A => X"0C2222C012488421884300000000000008CEFFF60F0000000CEEEEC01111111F",
            INIT_RAM_0B => X"137FFFFF0444E1008888888800000000888F888808CEFEC822222222088A7AC8",
            INIT_RAM_0C => X"111111115A5A5A5A00000000F00000000000000FFFFF00000000000000000000",
            INIT_RAM_0D => X"FF00000088880000000F8888FFFF0000888F88883333333300008CEF5A5A0000",
            INIT_RAM_0E => X"000000FF77777777000000000000000088888888888F0000000F8888888F0000",
            INIT_RAM_0F => X"FFFF000000000000000888880000FFFF00000000F1111111FFF0000000000FFF",
            INIT_RAM_10 => X"F3DD1FD3FFFF7FF1F1FF7FF1F7BDDDB7F3DFFFD3F3DD3DD3FDDD1DB7F1F395D3",
            INIT_RAM_11 => X"F7BDDDB7FDD95DDDFDDD559DF1FFFFFFFDB7F7BDF7BBBBB1F3777773FDDD1DDD",
            INIT_RAM_12 => X"FD955DDDF77BBDDDF3DDDDDDF7777771F3DD3FD3FDB73DD3F5B5DDB7FFFF3DD3",
            INIT_RAM_13 => X"FFF0FFFF7777537FF3BBBBB3F1FF3FF3F3FFFFF3F1FF7BD1F7773DDDFDDB7BDD",
            INIT_RAM_14 => X"FFFFFF7BF5B5F77FF99F7BDFF7353717FBB1B1BBFFFFFBBBF7FF7777FFFFFFFF",
            INIT_RAM_15 => X"FFFF7BDFF77FFFFFFFFF1FFFF77FFFFFFF77177FF7531357FFF777FFFB7FFF7B",
            INIT_RAM_16 => X"FFFF7BD1F3DD3FF3F7BDB7F1FBB1BB3BF3DD3DD3F1FF3DD3F1777777F3DD59D3",
            INIT_RAM_17 => X"FFFF3DD3FF73937FFFF1F1FFF17FFF71F77FF7FFFF7FF7FFF7BD1DD3F3DD3DD3",
            INIT_RAM_18 => X"FFFFFFFFFF0FFFFFFFFFFF0FFFFFF0FFFFFF0FFFFFFFFFFFF1300137FFF0FFFF",
            INIT_RAM_19 => X"FFFFFFF0FFFF7BDEEDB7FFFF0FFFFFFFFFFFF777FFFCB77777FFFFFFBBBBBBBB",
            INIT_RAM_1A => X"F3DDDD3FEDB77BDE77BCFFFFFFFFFFFFF7310009F0FFFFFFF311113FEEEEEEE0",
            INIT_RAM_1B => X"EC800000FBBB1EFF77777777FFFFFFFF77707777F7310137DDDDDDDDF7758537",
            INIT_RAM_1C => X"EEEEEEEEA5A5A5A5FFFFFFFF0FFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_1D => X"00FFFFFF7777FFFFFFF077770000FFFF77707777CCCCCCCCFFFF7310A5A5FFFF",
            INIT_RAM_1E => X"FFFFFF0088888888FFFFFFFFFFFFFFFF777777777770FFFFFFF077777770FFFF",
            INIT_RAM_1F => X"0000FFFFFFFFFFFFFFF77777FFFF0000FFFFFFFF0EEEEEEE000FFFFFFFFFF000",
            INIT_RAM_20 => X"C2A66A000000C02C0C0E2C000A626A220C202C000C222C000A4C48000E0C6A2C",
            INIT_RAM_21 => X"0C222C0002222C00099996000C8888880480840084444C040C88880802222C00",
            INIT_RAM_22 => X"06999100084222000A6222000C200C000C2C0E0000002C0022A66A0000C22C00",
            INIT_RAM_23 => X"000F00008888AC800C44444C0E00C00C0C00000C0E084E00C2A6220002484200",
            INIT_RAM_24 => X"000000840A4A08800660842008CAC8E8044E4E44000004440800888800000000",
            INIT_RAM_25 => X"00008420088000000000E000088000000088E88008ACECA80008880004800084",
            INIT_RAM_26 => X"0000842E0C22C00C0842480E044E44C40C22C22C0E00C22C0E8888880C22A62C",
            INIT_RAM_27 => X"0000C22C008C6C80000E0E000E80008E08800800008008000842E22C0C22C22C",
            INIT_RAM_28 => X"0C22E02C0000800E0E00800E084222480C20002C0C22C22C0222E248000F0000",
            INIT_RAM_29 => X"084222480226A2220222AA620E000000024808420844444E0C88888C0222E222",
            INIT_RAM_2A => X"026AA222088442220C2222220888888E0C22C02C0248C22C0A4A22480000C22C",
            INIT_RAM_2B => X"936C936C33CC33CC8888888800000000888F88880E00842E0888C22202248422",
            INIT_RAM_2C => X"111111115A5A5A5A00000000F00000000000000FFFFF00000000000000000000",
            INIT_RAM_2D => X"FF00000088880000000F8888FFFF0000888F888833333333C639C6395A5A0000",
            INIT_RAM_2E => X"000000FF77777777000000000000000088888888888F0000000F8888888F0000",
            INIT_RAM_2F => X"FFFF000000000000000888880000FFFF0000000000008421FFF0000000000FFF",
            INIT_RAM_30 => X"3D5995FFFFFF3FD3F3F1D3FFF59D95DDF3DFD3FFF3DDD3FFF5B3B7FFF1F395D3",
            INIT_RAM_31 => X"F3DDD3FFFDDDD3FFF66669FFF3777777FB7F7BFF7BBBB3FBF37777F7FDDDD3FF",
            INIT_RAM_32 => X"F9666EFFF7BDDDFFF59DDDFFF3DFF3FFF3D3F1FFFFFFD3FFDD5995FFFF3DD3FF",
            INIT_RAM_33 => X"FFF0FFFF7777537FF3BBBBB3F1FF3FF3F3FFFFF3F1F7B1FF3D59DDFFFDB7BDFF",
            INIT_RAM_34 => X"FFFFFF7BF5B5F77FF99F7BDFF7353717FBB1B1BBFFFFFBBBF7FF7777FFFFFFFF",
            INIT_RAM_35 => X"FFFF7BDFF77FFFFFFFFF1FFFF77FFFFFFF77177FF7531357FFF777FFFB7FFF7B",
            INIT_RAM_36 => X"FFFF7BD1F3DD3FF3F7BDB7F1FBB1BB3BF3DD3DD3F1FF3DD3F1777777F3DD59D3",
            INIT_RAM_37 => X"FFFF3DD3FF73937FFFF1F1FFF17FFF71F77FF7FFFF7FF7FFF7BD1DD3F3DD3DD3",
            INIT_RAM_38 => X"F3DD1FD3FFFF7FF1F1FF7FF1F7BDDDB7F3DFFFD3F3DD3DD3FDDD1DB7FFF0FFFF",
            INIT_RAM_39 => X"F7BDDDB7FDD95DDDFDDD559DF1FFFFFFFDB7F7BDF7BBBBB1F3777773FDDD1DDD",
            INIT_RAM_3A => X"FD955DDDF77BBDDDF3DDDDDDF7777771F3DD3FD3FDB73DD3F5B5DDB7FFFF3DD3",
            INIT_RAM_3B => X"6C936C93CC33CC3377777777FFFFFFFF77707777F1FF7BD1F7773DDDFDDB7BDD",
            INIT_RAM_3C => X"EEEEEEEEA5A5A5A5FFFFFFFF0FFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"00FFFFFF7777FFFFFFF077770000FFFF77707777CCCCCCCC39C639C6A5A5FFFF",
            INIT_RAM_3E => X"FFFFFF0088888888FFFFFFFFFFFFFFFF777777777770FFFFFFF077777770FFFF",
            INIT_RAM_3F => X"0000FFFFFFFFFFFFFFF77777FFFF0000FFFFFFFFFFFF7BDE000FFFFFFFFFF000"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 4,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0124442104447447074474470722222701244421072232270444742101245421",
            INIT_RAM_01 => X"0124442104444564044455640744444404447444034000000100000104447444",
            INIT_RAM_02 => X"0465544401122444034444440000000303403443044474470124442104447447",
            INIT_RAM_03 => X"0127210000002100030000030671311003222223074210070000122204421244",
            INIT_RAM_04 => X"0000010003443443042106600030121002272722000002220000000000000000",
            INIT_RAM_05 => X"0421000001100000000070001000000000003000002131200210001200011100",
            INIT_RAM_06 => X"0111004703447421034007470007210003401043074300430300021003465443",
            INIT_RAM_07 => X"0101004307100017000707000013631010000000000000000300344303443443",
            INIT_RAM_08 => X"2222222200F00000000000F000000F000000F0001111111103177310000F0000",
            INIT_RAM_09 => X"8888888F8421000000001248F8888888000E100000000000001E000000000000",
            INIT_RAM_0A => X"03444430842112480000000044444444001377730F000000037777300000000F",
            INIT_RAM_0B => X"0000137F01153000000000005A5A5A5A000F0000001373100000000000027210",
            INIT_RAM_0C => X"000000005A5A5A5A88888888F00000000000000FFFFF0000FFFFFFFF00000000",
            INIT_RAM_0D => X"FF000000000F0000000000000000000000000000000000008CEFFFFF5A5A0000",
            INIT_RAM_0E => X"000000FF00000000EEEEEEEECCCCCCCC000F0000000F0000000F000000000000",
            INIT_RAM_0F => X"0000FFFF0000FFFF000F000000000000FFFF0000F0000000FFF0000000000FFF",
            INIT_RAM_10 => X"FEDBBBDEFBBB8BB8F8BB8BB8F8DDDDD8FEDBBBDEF8DDCDD8FBBB8BDEFEDBABDE",
            INIT_RAM_11 => X"FEDBBBDEFBBBBA9BFBBBAA9BF8BBBBBBFBBB8BBBFCBFFFFFFEFFFFFEFBBB8BBB",
            INIT_RAM_12 => X"FB9AABBBFEEDDBBBFCBBBBBBFFFFFFFCFCBFCBBCFBBB8BB8FEDBBBDEFBBB8BB8",
            INIT_RAM_13 => X"FED8DEFFFFFFDEFFFCFFFFFCF98ECEEFFCDDDDDCF8BDEFF8FFFFEDDDFBBDEDBB",
            INIT_RAM_14 => X"FFFFFEFFFCBBCBBCFBDEF99FFFCFEDEFFDD8D8DDFFFFFDDDFFFFFFFFFFFFFFFF",
            INIT_RAM_15 => X"FBDEFFFFFEEFFFFFFFFF8FFFEFFFFFFFFFFFCFFFFFDECEDFFDEFFFEDFFFEEEFF",
            INIT_RAM_16 => X"FEEEFFB8FCBB8BDEFCBFF8B8FFF8DEFFFCBFEFBCF8BCFFBCFCFFFDEFFCB9ABBC",
            INIT_RAM_17 => X"FEFEFFBCF8EFFFE8FFF8F8FFFFEC9CEFEFFFFFFFFFFFFFFFFCFFCBBCFCBBCBBC",
            INIT_RAM_18 => X"DDDDDDDDFF0FFFFFFFFFFF0FFFFFF0FFFFFF0FFFEEEEEEEEFCE88CEFFFF0FFFF",
            INIT_RAM_19 => X"777777707BDEFFFFFFFFEDB707777777FFF1EFFFFFFFFFFFFFE1FFFFFFFFFFFF",
            INIT_RAM_1A => X"FCBBBBCF7BDEEDB7FFFFFFFFBBBBBBBBFFEC888CF0FFFFFFFC8888CFFFFFFFF0",
            INIT_RAM_1B => X"FFFFEC80FEEACFFFFFFFFFFFA5A5A5A5FFF0FFFFFFEC8CEFFFFFFFFFFFFD8DEF",
            INIT_RAM_1C => X"FFFFFFFFA5A5A5A5777777770FFFFFFFFFFFFFF00000FFFF00000000FFFFFFFF",
            INIT_RAM_1D => X"00FFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF73100000A5A5FFFF",
            INIT_RAM_1E => X"FFFFFF00FFFFFFFF1111111133333333FFF0FFFFFFF0FFFFFFF0FFFFFFFFFFFF",
            INIT_RAM_1F => X"FFFF0000FFFF0000FFF0FFFFFFFFFFFF0000FFFF0FFFFFFF000FFFFFFFFFF000",
            INIT_RAM_20 => X"3034430001117110034743000344430003444300056465440343030001245421",
            INIT_RAM_21 => X"0344430004446500044447000100000104654444340000000100010004446544",
            INIT_RAM_22 => X"0344440001244400034444000011171107034300044465000034430044566500",
            INIT_RAM_23 => X"0127210000002100030000030671311003222223072107003034440004212400",
            INIT_RAM_24 => X"0000010003443443042106600030121002272722000002220000000000000000",
            INIT_RAM_25 => X"0421000001100000000070001000000000003000002131200210001200011100",
            INIT_RAM_26 => X"0111004703447421034007470007210003401043074300430300021003465443",
            INIT_RAM_27 => X"0101004307100017000707000013631010000000000000000300344303443443",
            INIT_RAM_28 => X"01244421044474470744744707222227012444210722322704447421000F0000",
            INIT_RAM_29 => X"0124442104444564044455640744444404447444034000000100000104447444",
            INIT_RAM_2A => X"0465544401122444034444440000000303403443044474470124442104447447",
            INIT_RAM_2B => X"936C936C33CC33CC000000005A5A5A5A000F0000074210070000122204421244",
            INIT_RAM_2C => X"000000005A5A5A5A88888888F00000000000000FFFFF0000FFFFFFFF00000000",
            INIT_RAM_2D => X"FF000000000F000000000000000000000000000000000000C639C6395A5A0000",
            INIT_RAM_2E => X"000000FF00000000EEEEEEEECCCCCCCC000F0000000F0000000F000000000000",
            INIT_RAM_2F => X"0000FFFF0000FFFF000F000000000000FFFF000004654400FFF0000000000FFF",
            INIT_RAM_30 => X"CFCBBCFFFEEE8EEFFCB8BCFFFCBBBCFFFCBBBCFFFA9B9ABBFCBCFCFFFEDBABDE",
            INIT_RAM_31 => X"FCBBBCFFFBBB9AFFFBBBB8FFFEFFFFFEFB9ABBBBCBFFFFFFFEFFFEFFFBBB9ABB",
            INIT_RAM_32 => X"FCBBBBFFFEDBBBFFFCBBBBFFFFEEE8EEF8FCBCFFFBBB9AFFFFCBBCFFBBA99AFF",
            INIT_RAM_33 => X"FED8DEFFFFFFDEFFFCFFFFFCF98ECEEFFCDDDDDCF8DEF8FFCFCBBBFFFBDEDBFF",
            INIT_RAM_34 => X"FFFFFEFFFCBBCBBCFBDEF99FFFCFEDEFFDD8D8DDFFFFFDDDFFFFFFFFFFFFFFFF",
            INIT_RAM_35 => X"FBDEFFFFFEEFFFFFFFFF8FFFEFFFFFFFFFFFCFFFFFDECEDFFDEFFFEDFFFEEEFF",
            INIT_RAM_36 => X"FEEEFFB8FCBB8BDEFCBFF8B8FFF8DEFFFCBFEFBCF8BCFFBCFCFFFDEFFCB9ABBC",
            INIT_RAM_37 => X"FEFEFFBCF8EFFFE8FFF8F8FFFFEC9CEFEFFFFFFFFFFFFFFFFCFFCBBCFCBBCBBC",
            INIT_RAM_38 => X"FEDBBBDEFBBB8BB8F8BB8BB8F8DDDDD8FEDBBBDEF8DDCDD8FBBB8BDEFFF0FFFF",
            INIT_RAM_39 => X"FEDBBBDEFBBBBA9BFBBBAA9BF8BBBBBBFBBB8BBBFCBFFFFFFEFFFFFEFBBB8BBB",
            INIT_RAM_3A => X"FB9AABBBFEEDDBBBFCBBBBBBFFFFFFFCFCBFCBBCFBBB8BB8FEDBBBDEFBBB8BB8",
            INIT_RAM_3B => X"6C936C93CC33CC33FFFFFFFFA5A5A5A5FFF0FFFFF8BDEFF8FFFFEDDDFBBDEDBB",
            INIT_RAM_3C => X"FFFFFFFFA5A5A5A5777777770FFFFFFFFFFFFFF00000FFFF00000000FFFFFFFF",
            INIT_RAM_3D => X"00FFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF39C639C6A5A5FFFF",
            INIT_RAM_3E => X"FFFFFF00FFFFFFFF1111111133333333FFF0FFFFFFF0FFFFFFF0FFFFFFFFFFFF",
            INIT_RAM_3F => X"FFFF0000FFFF0000FFF0FFFFFFFFFFFF0000FFFFFB9ABBFF000FFFFFFFFFF000"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_1_AD_i
        );

end Behavioral; --Gowin_pROM_char
